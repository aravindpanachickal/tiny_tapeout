magic
tech sky130A
timestamp 1713328612
<< nwell >>
rect -56 -71 56 71
<< pmos >>
rect -9 -40 9 40
<< pdiff >>
rect -38 34 -9 40
rect -38 -34 -32 34
rect -15 -34 -9 34
rect -38 -40 -9 -34
rect 9 34 38 40
rect 9 -34 15 34
rect 32 -34 38 34
rect 9 -40 38 -34
<< pdiffc >>
rect -32 -34 -15 34
rect 15 -34 32 34
<< poly >>
rect -9 40 9 53
rect -9 -53 9 -40
<< locali >>
rect -32 34 -15 42
rect -32 -42 -15 -34
rect 15 34 32 42
rect 15 -42 32 -34
<< viali >>
rect -32 -34 -15 34
rect 15 -34 32 34
<< metal1 >>
rect -35 34 -12 40
rect -35 -34 -32 34
rect -15 -34 -12 34
rect -35 -40 -12 -34
rect 12 34 35 40
rect 12 -34 15 34
rect 32 -34 35 34
rect 12 -40 35 -34
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.8 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
