magic
tech sky130A
<<<<<<< HEAD
timestamp 1713437673
=======
timestamp 1713438817
>>>>>>> d91cb2988effe7e4f0e56e7a27fb6a110da9f303
<< error_p >>
rect -56 -193 56 193
<< nwell >>
rect -56 -193 56 193
<< pmos >>
rect -9 -162 9 162
<< pdiff >>
rect -38 156 -9 162
rect -38 -156 -32 156
rect -15 -156 -9 156
rect -38 -162 -9 -156
rect 9 156 38 162
rect 9 -156 15 156
rect 32 -156 38 156
rect 9 -162 38 -156
<< pdiffc >>
rect -32 -156 -15 156
rect 15 -156 32 156
<< poly >>
rect -9 162 9 175
rect -9 -175 9 -162
<< locali >>
rect -32 156 -15 164
rect -32 -164 -15 -156
rect 15 156 32 164
rect 15 -164 32 -156
<< viali >>
rect -32 -156 -15 156
rect 15 -156 32 156
<< metal1 >>
rect -35 156 -12 162
rect -35 -156 -32 156
rect -15 -156 -12 156
rect -35 -162 -12 -156
rect 12 156 35 162
rect 12 -156 15 156
rect 32 -156 35 156
rect 12 -162 35 -156
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.24 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
