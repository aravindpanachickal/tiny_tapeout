magic
tech sky130A
magscale 1 2

<< nwell >>
rect -590 1930 2556 2520
rect 124 1893 299 1930
rect 1048 1889 2556 1930
rect 1048 1583 2553 1889

<< ndiff >>
rect -402 1574 -2 1600
rect 427 1499 728 1524
rect 2651 1509 2951 1535
rect 1396 1181 1696 1206
rect 1406 718 1706 744
rect 2161 721 2463 751
<< pdiff >>
rect -529 2122 121 2153
rect 349 2140 966 2154
rect 317 2126 966 2140
rect 1208 2125 1858 2153
rect 2132 2124 2372 2151
rect 2161 1668 2321 1699
rect 1226 1628 1874 1655
<< psubdiff >>
rect -402 1553 -2 1574
rect -402 1490 -340 1553
rect -60 1490 -2 1553
rect -402 1464 -2 1490
rect 427 1457 728 1499
rect 427 1396 446 1457
rect 705 1396 728 1457
rect 427 1344 728 1396
rect 2651 1480 2951 1509
rect 2651 1421 2680 1480
rect 2930 1421 2951 1480
rect 2651 1380 2951 1421
rect 1396 1150 1696 1181
rect 1396 1091 1422 1150
rect 1672 1091 1696 1150
rect 1396 1057 1696 1091
rect 1406 691 1706 718
rect 1406 632 1431 691
rect 1681 632 1706 691
rect 1406 590 1706 632
rect 2161 688 2463 721
rect 2161 629 2189 688
rect 2439 629 2463 688
rect 2161 590 2463 629
<< nsubdiff >>
rect -529 2371 121 2441
rect -529 2227 -414 2371
rect 4 2227 121 2371
rect -529 2153 121 2227
rect 317 2379 966 2439
rect 317 2235 432 2379
rect 850 2235 966 2379
rect 317 2154 966 2235
rect 317 2140 349 2154
rect 1208 2390 1858 2417
rect 1208 2246 1327 2390
rect 1745 2246 1858 2390
rect 1208 2153 1858 2246
rect 2132 2342 2372 2427
rect 2132 2248 2204 2342
rect 2308 2248 2372 2342
rect 2132 2151 2372 2248
rect 1226 1821 1874 1860
rect 1226 1677 1341 1821
rect 1759 1677 1874 1821
rect 1226 1655 1874 1677
rect 2161 1751 2321 1780
rect 2161 1716 2202 1751
rect 2281 1716 2321 1751
rect 2161 1699 2321 1716
<< psubdiffcont >>
rect -340 1490 -60 1553
rect 446 1396 705 1457
rect 2680 1421 2930 1480
rect 1422 1091 1672 1150
rect 1431 632 1681 691
rect 2189 629 2439 688
<< nsubdiffcont >>
rect -414 2227 4 2371
rect 432 2235 850 2379
rect 1327 2246 1745 2390
rect 2204 2248 2308 2342
rect 1341 1677 1759 1821
rect 2202 1716 2281 1751
<< poly >>
rect 139 2034 300 2071
rect 1085 2070 1152 2093
rect 2439 2073 2505 2088
rect 1085 2069 1199 2070
rect 2439 2069 2455 2073
rect 1085 2035 1102 2069
rect 1136 2035 1199 2069
rect 1085 2034 1199 2035
rect 2395 2039 2455 2069
rect 2489 2039 2505 2073
rect 192 1961 233 2034
rect 1085 2008 1152 2034
rect 2395 2033 2505 2039
rect 2439 2020 2505 2033
rect 180 1950 247 1961
rect 180 1916 196 1950
rect 231 1916 247 1950
rect 180 1906 247 1916
rect -511 1693 -451 1715
rect -511 1654 -499 1693
rect -465 1657 -410 1693
rect -465 1654 -451 1657
rect -511 1636 -451 1654
rect 288 1618 380 1645
rect 288 1614 409 1618
rect 288 1580 316 1614
rect 351 1582 409 1614
rect 2059 1616 2122 1631
rect 2536 1628 2610 1654
rect 2059 1615 2141 1616
rect 351 1580 380 1582
rect 288 1549 380 1580
rect 1087 1572 1161 1591
rect 2059 1581 2074 1615
rect 2108 1581 2141 1615
rect 2059 1580 2141 1581
rect 2536 1594 2564 1628
rect 2598 1594 2630 1628
rect 2536 1592 2630 1594
rect 1087 1571 1213 1572
rect 1087 1537 1105 1571
rect 1139 1537 1213 1571
rect 2059 1564 2122 1580
rect 2536 1574 2610 1592
rect 1087 1536 1213 1537
rect 1087 1512 1161 1536
rect 1267 1300 1328 1316
rect 1267 1299 1386 1300
rect 1267 1265 1280 1299
rect 1314 1265 1386 1299
rect 1267 1264 1386 1265
rect 1267 1245 1328 1264
rect 1291 837 1359 856
rect 2067 840 2122 861
rect 1291 803 1306 837
rect 1340 803 1397 837
rect 1291 801 1397 803
rect 2067 806 2077 840
rect 2111 806 2156 840
rect 2067 804 2156 806
rect 1291 786 1359 801
rect 2067 785 2122 804
<< polycont >>
rect 1102 2035 1136 2069
rect 2455 2039 2489 2073
rect 196 1916 231 1950
rect -499 1654 -465 1693
rect 316 1580 351 1614
rect 2074 1581 2108 1615
rect 2564 1594 2598 1628
rect 1105 1537 1139 1571
rect 1280 1265 1314 1299
rect 1306 803 1340 837
rect 2077 806 2111 840
<< locali >>
rect -529 2745 121 2810
rect -529 2594 -289 2745
rect -122 2594 121 2745
rect -529 2371 121 2594
rect -529 2227 -414 2371
rect 4 2227 121 2371
rect -529 2115 121 2227
rect 316 2743 966 2810
rect 316 2592 566 2743
rect 733 2592 966 2743
rect 316 2379 966 2592
rect 316 2235 432 2379
rect 850 2235 966 2379
rect 316 2113 966 2235
rect 1208 2742 1858 2810
rect 1208 2591 1444 2742
rect 1611 2591 1858 2742
rect 1208 2390 1858 2591
rect 1208 2246 1327 2390
rect 1745 2246 1858 2390
rect 1208 2114 1858 2246
rect 2132 2738 2372 2810
rect 2132 2587 2173 2738
rect 2340 2587 2372 2738
rect 2132 2342 2372 2587
rect 2132 2248 2204 2342
rect 2308 2248 2372 2342
rect 2132 2109 2372 2248
rect 1085 2069 1152 2093
rect 1085 2035 1102 2069
rect 1136 2035 1152 2069
rect -389 1869 -13 2017
rect 180 1950 247 1961
rect 180 1916 196 1950
rect 231 1916 247 1950
rect 180 1906 247 1916
rect 192 1869 235 1906
rect -389 1832 235 1869
rect 549 1868 625 2013
rect 1085 2008 1152 2035
rect 2439 2075 2505 2088
rect 2564 2075 2606 2076
rect 2439 2073 2606 2075
rect 2439 2039 2455 2073
rect 2489 2041 2606 2073
rect 2489 2039 2505 2041
rect 2439 2020 2505 2039
rect 549 1865 989 1868
rect -511 1693 -451 1715
rect -389 1712 -13 1832
rect 549 1818 991 1865
rect -511 1691 -499 1693
rect -582 1655 -499 1691
rect -511 1654 -499 1655
rect -465 1654 -451 1693
rect 948 1664 991 1818
rect -511 1636 -451 1654
rect 288 1632 380 1645
rect -402 1553 -2 1611
rect -402 1490 -340 1553
rect -60 1490 -2 1553
rect 288 1566 300 1632
rect 370 1566 380 1632
rect 729 1630 992 1664
rect 288 1549 380 1566
rect -402 1464 -2 1490
rect -400 461 -2 1464
rect 427 1457 728 1560
rect 427 1396 446 1457
rect 705 1396 728 1457
rect 427 1344 728 1396
rect 948 1399 991 1630
rect 1105 1591 1139 2008
rect 1277 1932 1836 2019
rect 2227 1948 2261 2018
rect 1277 1898 2051 1932
rect 2226 1907 2261 1948
rect 1277 1860 1836 1898
rect 1226 1821 1874 1860
rect 1226 1677 1341 1821
rect 1759 1677 1874 1821
rect 2017 1781 2051 1898
rect 2213 1892 2278 1907
rect 2213 1850 2225 1892
rect 2265 1850 2278 1892
rect 2213 1839 2278 1850
rect 2017 1780 2319 1781
rect 2017 1751 2321 1780
rect 2564 1762 2606 2041
rect 2017 1747 2202 1751
rect 1226 1614 1874 1677
rect 2161 1716 2202 1747
rect 2281 1716 2321 1751
rect 2161 1658 2321 1716
rect 2430 1728 2606 1762
rect 2059 1615 2122 1631
rect 1086 1571 1161 1591
rect 1086 1537 1105 1571
rect 1139 1537 1161 1571
rect 2059 1581 2074 1615
rect 2108 1581 2122 1615
rect 2059 1564 2122 1581
rect 1086 1512 1161 1537
rect 1108 1399 1142 1512
rect 1402 1434 1678 1520
rect 1402 1399 1843 1434
rect 948 1363 1143 1399
rect 951 1362 1143 1363
rect -400 380 -341 461
rect -68 380 -2 461
rect -400 342 -2 380
rect 438 468 710 1344
rect 1108 1308 1142 1362
rect 438 390 498 468
rect 652 390 710 468
rect 438 342 710 390
rect 1107 1300 1142 1308
rect 1267 1300 1328 1316
rect 1402 1313 1678 1399
rect 1809 1326 1843 1399
rect 1107 1299 1328 1300
rect 1107 1266 1280 1299
rect 1107 837 1142 1266
rect 1267 1265 1280 1266
rect 1314 1265 1328 1299
rect 1809 1288 1844 1326
rect 1267 1245 1328 1265
rect 1396 1150 1696 1247
rect 1810 1214 1844 1288
rect 2073 1214 2109 1564
rect 2224 1403 2258 1545
rect 2210 1383 2279 1403
rect 2210 1348 2226 1383
rect 2261 1348 2279 1383
rect 2210 1333 2279 1348
rect 2430 1214 2476 1728
rect 2564 1654 2606 1728
rect 2739 1776 2828 1795
rect 2739 1739 2765 1776
rect 2807 1739 2828 1776
rect 2739 1721 2828 1739
rect 2760 1674 2802 1721
rect 2536 1628 2610 1654
rect 2647 1641 2802 1674
rect 2647 1640 2783 1641
rect 2536 1594 2564 1628
rect 2598 1594 2610 1628
rect 2536 1574 2610 1594
rect 2651 1480 2951 1577
rect 2651 1421 2680 1480
rect 2930 1421 2951 1480
rect 2651 1380 2951 1421
rect 1810 1180 2476 1214
rect 1396 1091 1422 1150
rect 1672 1091 1696 1150
rect 1396 1057 1696 1091
rect 1425 997 1668 1057
rect 1425 995 1949 997
rect 1425 961 1950 995
rect 1425 860 1668 961
rect 1291 837 1359 856
rect 1107 803 1306 837
rect 1340 803 1359 837
rect 1107 802 1359 803
rect 1107 29 1150 802
rect 1291 786 1359 802
rect 1406 691 1706 783
rect 1406 632 1431 691
rect 1681 632 1706 691
rect 1406 590 1706 632
rect 1909 664 1950 961
rect 2073 861 2111 1180
rect 2153 1179 2437 1180
rect 2266 1006 2355 1019
rect 2266 961 2289 1006
rect 2328 961 2355 1006
rect 2266 945 2355 961
rect 2287 861 2331 945
rect 2067 840 2122 861
rect 2067 806 2077 840
rect 2111 806 2122 840
rect 2067 785 2122 806
rect 2161 688 2463 789
rect 2161 664 2189 688
rect 1909 629 2189 664
rect 2439 629 2463 688
rect 1909 627 2463 629
rect 2161 590 2463 627
rect 1408 464 1705 590
rect 1408 380 1439 464
rect 1669 380 1705 464
rect 1408 342 1705 380
rect 2652 474 2950 1380
rect 2652 383 2737 474
rect 2877 383 2950 474
rect 2652 342 2950 383
rect -560 -15 -202 21
rect -560 -170 -490 -15
rect -269 -170 -202 -15
rect -560 -209 -202 -170
rect 943 -8 1276 29
rect 943 -175 1006 -8
rect 1209 -175 1276 -8
rect 943 -205 1276 -175
rect -519 -466 -236 -209
rect -519 -749 3149 -466
rect -5669 -879 -5029 -750
rect -5669 -1178 -5506 -879
rect -5154 -901 -5029 -879
rect 2866 -901 3149 -749
rect -5154 -1178 -4755 -901
rect -5669 -1183 -4755 -1178
rect -5669 -1308 -5029 -1183
<< viali >>
rect -289 2594 -122 2745
rect 566 2592 733 2743
rect 1444 2591 1611 2742
rect 2173 2587 2340 2738
rect 300 1614 370 1632
rect 300 1580 316 1614
rect 316 1580 351 1614
rect 351 1580 370 1614
rect 300 1566 370 1580
rect 2225 1850 2265 1892
rect -341 380 -68 461
rect 498 390 652 468
rect 2226 1348 2261 1383
rect 2765 1739 2807 1776
rect 2289 961 2328 1006
rect 1439 380 1669 464
rect 2737 383 2877 474
rect -490 -170 -269 -15
rect 1006 -175 1209 -8
rect -5506 -1178 -5154 -879
<< metal1 >>
rect -590 2745 2547 2810
rect -590 2594 -289 2745
rect -122 2743 2547 2745
rect -122 2594 566 2743
rect -590 2592 566 2594
rect 733 2742 2547 2743
rect 733 2592 1444 2742
rect -590 2591 1444 2592
rect 1611 2738 2547 2742
rect 1611 2591 2173 2738
rect -590 2587 2173 2591
rect 2340 2587 2547 2738
rect -590 2530 2547 2587
rect 315 2384 3085 2421
rect 316 2213 349 2384
rect 317 1662 349 2213
rect 2213 1892 2278 1907
rect 2213 1850 2225 1892
rect 2265 1886 2278 1892
rect 3051 1886 3085 2384
rect 2265 1858 3342 1886
rect 2265 1857 3085 1858
rect 3155 1857 3342 1858
rect 2265 1850 2278 1857
rect 2213 1839 2278 1850
rect 2770 1795 2798 1857
rect 2739 1776 2828 1795
rect 2739 1739 2765 1776
rect 2807 1739 2828 1776
rect 2739 1721 2828 1739
rect 272 1632 395 1662
rect 272 1566 300 1632
rect 370 1566 395 1632
rect 272 1529 395 1566
rect 317 1528 360 1529
rect 2210 1383 2279 1403
rect 2210 1348 2226 1383
rect 2261 1348 2279 1383
rect 2210 1333 2279 1348
rect 2221 1296 2269 1333
rect 1968 1248 2269 1296
rect 1968 498 2016 1248
rect 2266 1008 2355 1019
rect 2266 1006 3194 1008
rect 2266 961 2289 1006
rect 2328 967 3194 1006
rect 2328 961 2355 967
rect 2266 945 2355 961
rect -560 474 2952 498
rect -560 468 2737 474
rect -560 461 498 468
rect -560 380 -341 461
rect -68 390 498 461
rect 652 464 2737 468
rect 652 390 1439 464
rect -68 380 1439 390
rect 1669 383 2737 464
rect 2877 383 2952 474
rect 1669 380 2952 383
rect -560 342 2952 380
rect -560 -15 -202 342
rect -560 -170 -490 -15
rect -269 -170 -202 -15
rect -560 -209 -202 -170
rect 943 -8 1276 29
rect 943 -175 1006 -8
rect 1209 -175 1276 -8
rect 943 -205 1276 -175
rect -5669 -879 -5029 -750
rect -5669 -1178 -5506 -879
rect -5154 -1178 -5029 -879
rect -5669 -1308 -5029 -1178
<< via1 >>
rect -490 -170 -269 -15
rect 1006 -175 1209 -8
rect -5506 -1178 -5154 -879
<< metal2 >>
rect -560 -15 -202 21
rect -560 -170 -490 -15
rect -269 -170 -202 -15
rect -560 -209 -202 -170
rect 943 -8 1276 29
rect 943 -175 1006 -8
rect 1209 -175 1276 -8
rect 943 -205 1276 -175
rect -5669 -879 -5029 -750
rect -5669 -1178 -5506 -879
rect -5154 -1178 -5029 -879
rect -5669 -1308 -5029 -1178
<< via2 >>
rect -490 -170 -269 -15
rect 1006 -175 1209 -8
rect -5506 -1178 -5154 -879
<< metal3 >>
rect -542 -15 -202 21
rect -542 -67 -490 -15
rect -785 -150 -490 -67
rect -542 -170 -490 -150
rect -269 -170 -202 -15
rect -542 -209 -202 -170
rect 943 -8 1276 29
rect 943 -175 1006 -8
rect 1209 -175 1276 -8
rect 943 -205 1276 -175
rect -5669 -879 -5029 -750
rect -5669 -1178 -5506 -879
rect -5154 -1178 -5029 -879
rect -5669 -1308 -5029 -1178
<< via3 >>
rect 1006 -175 1209 -8
rect -5506 -1178 -5154 -879
<< metal4 >>
rect 943 -8 1276 29
rect 943 -175 1006 -8
rect 1209 -175 1276 -8
rect 943 -205 1276 -175
rect -5510 -750 -5227 -513
rect -1347 -693 -1155 -512
rect 1006 -693 1210 -205
rect -1347 -696 1210 -693
rect -5669 -879 -5029 -750
rect -1347 -856 1203 -696
rect -5669 -1178 -5506 -879
rect -5154 -1178 -5029 -879
rect -5669 -1308 -5029 -1178
use sky130_fd_pr__cap_mim_m3_1_MWYMHE  sky130_fd_pr__cap_mim_m3_1_MWYMHE_0

transform 0 -1 -779 1 0 -1042
box -141 -3976 141 3976
<< end >>
