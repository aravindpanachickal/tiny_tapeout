magic
tech sky130A
timestamp 1713328612
<< nmos >>
rect -9 -100 9 100
<< ndiff >>
rect -38 94 -9 100
rect -38 -94 -32 94
rect -15 -94 -9 94
rect -38 -100 -9 -94
rect 9 94 38 100
rect 9 -94 15 94
rect 32 -94 38 94
rect 9 -100 38 -94
<< ndiffc >>
rect -32 -94 -15 94
rect 15 -94 32 94
<< poly >>
rect -9 100 9 113
rect -9 -113 9 -100
<< locali >>
rect -32 94 -15 102
rect -32 -102 -15 -94
rect 15 94 32 102
rect 15 -102 32 -94
<< viali >>
rect -32 -94 -15 94
rect 15 -94 32 94
<< metal1 >>
rect -35 94 -12 100
rect -35 -94 -32 94
rect -15 -94 -12 94
rect -35 -100 -12 -94
rect 12 94 35 100
rect 12 -94 15 94
rect 32 -94 35 94
rect 12 -100 35 -94
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
