magic
tech sky130A

<< error_p >>
rect -38 -75 -9 75
rect 9 -75 38 75
<< nmos >>
rect -9 -75 9 75
<< ndiff >>
rect -38 69 -9 75
rect -38 -69 -32 69
rect -15 -69 -9 69
rect -38 -75 -9 -69
rect 9 69 38 75
rect 9 -69 15 69
rect 32 -69 38 69
rect 9 -75 38 -69
<< ndiffc >>
rect -32 -69 -15 69
rect 15 -69 32 69
<< poly >>
rect -9 75 9 88
rect -9 -88 9 -75
<< locali >>
rect -32 69 -15 77
rect -32 -77 -15 -69
rect 15 69 32 77
rect 15 -77 32 -69
<< viali >>
rect -32 -69 -15 69
rect 15 -69 32 69
<< metal1 >>
rect -35 69 -12 75
rect -35 -69 -32 69
rect -15 -69 -12 69
rect -35 -75 -12 -69
rect 12 69 35 75
rect 12 -69 15 69
rect 32 -69 35 69
rect 12 -75 35 -69
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.5 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
