magic
tech sky130A
magscale 1 2
timestamp 1713328612
<< pwell >>
rect -307 -4142 307 4142
<< psubdiff >>
rect -271 4072 -175 4106
rect 175 4072 271 4106
rect -271 4010 -237 4072
rect 237 4010 271 4072
rect -271 -4072 -237 -4010
rect 237 -4072 271 -4010
rect -271 -4106 -175 -4072
rect 175 -4106 271 -4072
<< psubdiffcont >>
rect -175 4072 175 4106
rect -271 -4010 -237 4010
rect 237 -4010 271 4010
rect -175 -4106 175 -4072
<< xpolycontact >>
rect -141 3544 141 3976
rect -141 -3976 141 -3544
<< xpolyres >>
rect -141 -3544 141 3544
<< locali >>
rect -271 4072 -175 4106
rect 175 4072 271 4106
rect -271 4010 -237 4072
rect 237 4010 271 4072
rect -271 -4072 -237 -4010
rect 237 -4072 271 -4010
rect -271 -4106 -175 -4072
rect 175 -4106 271 -4072
<< viali >>
rect -125 3561 125 3958
rect -125 -3958 125 -3561
<< metal1 >>
rect -131 3958 131 3970
rect -131 3561 -125 3958
rect 125 3561 131 3958
rect -131 3549 131 3561
rect -131 -3561 131 -3549
rect -131 -3958 -125 -3561
rect 125 -3958 131 -3561
rect -131 -3970 131 -3958
<< properties >>
string FIXED_BBOX -254 -4089 254 4089
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 35.441 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 50.537k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
