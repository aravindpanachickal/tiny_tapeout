magic
tech sky130A
magscale 1 2
timestamp 1713435522
<< nwell >>
rect 18679 4227 19528 4270
<< poly >>
rect 17016 4436 17147 4515
<< locali >>
rect 17016 4502 17147 4515
rect 17016 4449 17063 4502
rect 17134 4449 17147 4502
rect 17016 4436 17147 4449
rect 20354 4441 20358 4474
rect 20245 4440 20400 4441
<< viali >>
rect 17063 4449 17134 4502
<< metal1 >>
rect 842 5624 1435 5755
rect 842 5344 977 5624
rect 1312 5610 1435 5624
rect 1312 5344 17286 5610
rect 842 5330 17286 5344
rect 842 5245 1435 5330
rect 20911 4657 31384 4686
rect 17016 4502 17147 4515
rect 17016 4449 17063 4502
rect 17134 4449 17147 4502
rect 17016 4436 17147 4449
rect 20745 3767 26978 3808
rect 10328 3298 10537 3343
rect 10328 3286 17167 3298
rect 10328 3147 10376 3286
rect 10495 3147 17167 3286
rect 10328 3142 17167 3147
rect 10328 3095 10537 3142
rect 26937 460 26978 3767
rect 26880 438 27036 460
rect 31355 456 31383 4657
rect 26880 360 26920 438
rect 27002 360 27036 438
rect 26880 330 27036 360
rect 31298 428 31452 456
rect 31298 356 31330 428
rect 31424 356 31452 428
rect 31298 324 31452 356
<< via1 >>
rect 977 5344 1312 5624
rect 17063 4449 17134 4502
rect 10376 3147 10495 3286
rect 26920 360 27002 438
rect 31330 356 31424 428
<< metal2 >>
rect 842 5624 1435 5755
rect 842 5344 977 5624
rect 1312 5344 1435 5624
rect 842 5245 1435 5344
rect 17016 4502 17147 4515
rect 17016 4449 17063 4502
rect 17134 4449 17147 4502
rect 17016 4436 17147 4449
rect 10328 3286 10537 3343
rect 10328 3147 10376 3286
rect 10495 3147 10537 3286
rect 10328 3095 10537 3147
rect 17042 2994 17090 4436
rect 17042 2946 22584 2994
rect 22536 660 22584 2946
rect 22480 637 22600 660
rect 22480 570 22513 637
rect 22577 570 22600 637
rect 22480 544 22600 570
rect 26880 438 27036 460
rect 26880 360 26920 438
rect 27002 360 27036 438
rect 26880 330 27036 360
rect 31298 428 31452 456
rect 31298 356 31330 428
rect 31424 356 31452 428
rect 31298 324 31452 356
<< via2 >>
rect 977 5344 1312 5624
rect 10376 3147 10495 3286
rect 22513 570 22577 637
rect 26920 360 27002 438
rect 31330 356 31424 428
<< metal3 >>
rect 842 5624 1435 5755
rect 842 5344 977 5624
rect 1312 5344 1435 5624
rect 842 5245 1435 5344
rect 10328 3286 10537 3343
rect 10328 3147 10376 3286
rect 10495 3147 10537 3286
rect 10328 3095 10537 3147
rect 22480 637 22600 660
rect 22480 570 22513 637
rect 22577 570 22600 637
rect 22480 544 22600 570
rect 26880 438 27036 460
rect 26880 360 26920 438
rect 27002 360 27036 438
rect 26880 330 27036 360
rect 31298 428 31452 456
rect 31298 356 31330 428
rect 31424 356 31452 428
rect 31298 324 31452 356
<< via3 >>
rect 977 5344 1312 5624
rect 10376 3147 10495 3286
rect 22513 570 22577 637
rect 26920 360 27002 438
rect 31330 356 31424 428
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 5608 500 44152
rect 842 5624 1435 5755
rect 842 5608 977 5624
rect 200 5344 977 5608
rect 1312 5344 1435 5624
rect 200 5331 1435 5344
rect 200 1000 500 5331
rect 842 5245 1435 5331
rect 9800 3298 10100 44152
rect 10328 3298 10537 3343
rect 9800 3286 10537 3298
rect 9800 3147 10376 3286
rect 10495 3147 10537 3286
rect 9800 3141 10537 3147
rect 9800 1000 10100 3141
rect 10328 3095 10537 3141
rect 22480 637 22600 660
rect 22480 570 22513 637
rect 22577 570 22600 637
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 570
rect 26880 438 27036 460
rect 26880 360 26920 438
rect 27002 360 27036 438
rect 26880 330 27036 360
rect 31298 428 31452 456
rect 31298 356 31330 428
rect 31424 356 31452 428
rect 26896 0 27016 330
rect 31298 324 31452 356
rect 31312 0 31432 324
use leakylayout  leakylayout_0
timestamp 1713435522
transform 1 0 17598 0 1 2800
box -6357 -1308 3342 3486
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
