VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_analog_example
  CLASS BLOCK ;
  FOREIGN tt_um_analog_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.976400 ;
    ANTENNADIFFAREA 28.198374 ;
    PORT
      LAYER nwell ;
        RECT 88.560 23.770 104.290 26.720 ;
        RECT 92.130 23.585 93.005 23.770 ;
        RECT 96.915 23.565 104.290 23.770 ;
        RECT 96.915 22.035 104.275 23.565 ;
        RECT 96.915 21.555 104.270 22.035 ;
        RECT 96.915 21.360 104.250 21.555 ;
        RECT 96.915 21.330 102.620 21.360 ;
        RECT 101.125 21.295 102.620 21.330 ;
        RECT 101.125 21.270 102.555 21.295 ;
      LAYER li1 ;
        RECT 88.865 24.700 92.115 28.170 ;
        RECT 93.090 24.705 96.340 28.170 ;
        RECT 88.850 24.530 92.130 24.700 ;
        RECT 93.080 24.535 96.360 24.705 ;
        RECT 97.550 24.700 100.800 28.170 ;
        RECT 93.080 24.065 96.360 24.235 ;
        RECT 96.935 24.160 97.270 24.585 ;
        RECT 97.530 24.530 100.810 24.700 ;
        RECT 102.170 24.695 103.370 28.170 ;
        RECT 102.150 24.525 103.390 24.695 ;
        RECT 94.255 23.460 94.635 24.065 ;
        RECT 94.255 23.445 96.455 23.460 ;
        RECT 94.255 23.210 96.465 23.445 ;
        RECT 96.250 22.440 96.465 23.210 ;
        RECT 92.950 21.865 93.410 22.345 ;
        RECT 93.630 22.270 96.470 22.440 ;
        RECT 96.250 21.115 96.465 22.270 ;
        RECT 97.035 22.075 97.205 24.160 ;
        RECT 97.530 24.060 100.810 24.230 ;
        RECT 97.895 23.780 100.690 24.060 ;
        RECT 102.150 24.055 103.390 24.225 ;
        RECT 102.645 23.860 102.815 24.055 ;
        RECT 97.895 23.610 101.765 23.780 ;
        RECT 102.640 23.655 102.815 23.860 ;
        RECT 97.895 23.420 100.690 23.610 ;
        RECT 97.640 22.210 100.880 23.420 ;
        RECT 101.595 23.025 101.765 23.610 ;
        RECT 102.575 23.315 102.900 23.655 ;
        RECT 101.595 23.020 103.105 23.025 ;
        RECT 101.595 22.855 103.115 23.020 ;
        RECT 102.315 22.430 103.115 22.855 ;
        RECT 105.205 22.725 105.650 23.095 ;
        RECT 105.310 22.490 105.520 22.725 ;
        RECT 102.295 22.260 103.135 22.430 ;
        RECT 104.745 22.320 106.285 22.490 ;
        RECT 96.940 21.680 97.315 22.075 ;
        RECT 97.620 22.040 100.900 22.210 ;
        RECT 97.050 21.115 97.220 21.680 ;
        RECT 96.250 20.935 97.225 21.115 ;
        RECT 96.265 20.930 97.225 20.935 ;
        RECT 97.050 20.685 97.220 20.930 ;
        RECT 97.845 20.685 98.150 20.765 ;
        RECT 97.050 20.660 98.150 20.685 ;
        RECT 97.045 20.515 98.150 20.660 ;
        RECT 97.045 18.305 97.220 20.515 ;
        RECT 97.845 20.410 98.150 20.515 ;
        RECT 97.965 18.305 98.305 18.400 ;
        RECT 97.045 18.130 98.305 18.305 ;
        RECT 97.045 14.265 97.260 18.130 ;
        RECT 97.965 18.050 98.305 18.130 ;
        RECT 96.225 13.095 97.890 14.265 ;
        RECT 63.165 9.615 66.365 10.370 ;
        RECT 63.165 8.205 69.895 9.615 ;
        RECT 63.165 7.580 66.365 8.205 ;
      LAYER mcon ;
        RECT 90.065 27.090 90.900 27.845 ;
        RECT 94.340 27.080 95.175 27.835 ;
        RECT 98.730 27.075 99.565 27.830 ;
        RECT 88.930 24.530 92.050 24.700 ;
        RECT 93.160 24.535 96.280 24.705 ;
        RECT 102.375 27.055 103.210 27.810 ;
        RECT 93.160 24.065 96.280 24.235 ;
        RECT 97.610 24.530 100.730 24.700 ;
        RECT 102.230 24.525 103.310 24.695 ;
        RECT 93.010 21.950 93.360 22.280 ;
        RECT 93.710 22.270 95.090 22.440 ;
        RECT 97.610 24.060 100.730 24.230 ;
        RECT 102.230 24.055 103.310 24.225 ;
        RECT 102.635 23.370 102.835 23.580 ;
        RECT 105.335 22.815 105.545 23.000 ;
        RECT 102.375 22.260 103.055 22.430 ;
        RECT 104.825 22.320 106.205 22.490 ;
        RECT 97.700 22.040 100.820 22.210 ;
        RECT 96.540 13.245 97.555 14.080 ;
        RECT 63.980 8.230 65.740 9.725 ;
        RECT 67.825 8.285 69.810 9.535 ;
      LAYER met1 ;
        RECT 5.860 28.170 9.370 29.165 ;
        RECT 88.295 28.170 88.815 28.175 ;
        RECT 5.860 26.770 104.245 28.170 ;
        RECT 5.860 25.430 9.370 26.770 ;
        RECT 88.295 26.760 88.815 26.770 ;
        RECT 93.085 26.040 106.935 26.225 ;
        RECT 93.090 25.185 93.255 26.040 ;
        RECT 93.095 24.735 93.255 25.185 ;
        RECT 88.870 24.500 92.110 24.730 ;
        RECT 93.095 24.505 96.340 24.735 ;
        RECT 93.095 24.265 93.255 24.505 ;
        RECT 97.550 24.500 100.790 24.730 ;
        RECT 102.170 24.495 103.370 24.725 ;
        RECT 93.095 24.035 96.340 24.265 ;
        RECT 93.095 22.430 93.255 24.035 ;
        RECT 97.550 24.030 100.790 24.260 ;
        RECT 102.170 24.025 103.370 24.255 ;
        RECT 102.575 23.550 102.900 23.655 ;
        RECT 106.765 23.550 106.935 26.040 ;
        RECT 102.575 23.410 157.020 23.550 ;
        RECT 102.575 23.405 106.935 23.410 ;
        RECT 107.285 23.405 157.020 23.410 ;
        RECT 102.575 23.315 102.900 23.405 ;
        RECT 105.360 23.095 105.500 23.405 ;
        RECT 107.690 23.400 157.020 23.405 ;
        RECT 105.205 22.725 105.650 23.095 ;
        RECT 92.870 21.765 93.485 22.430 ;
        RECT 93.650 22.240 95.150 22.470 ;
        RECT 97.640 22.010 100.880 22.240 ;
        RECT 102.315 22.230 103.115 22.460 ;
        RECT 104.765 22.290 106.265 22.520 ;
        RECT 93.095 21.760 93.310 21.765 ;
        RECT 96.225 13.095 97.890 14.265 ;
        RECT 63.165 7.580 66.365 10.370 ;
        RECT 67.765 8.255 69.870 9.565 ;
        RECT 156.730 2.060 157.020 23.400 ;
        RECT 156.420 1.320 157.310 2.060 ;
      LAYER via ;
        RECT 6.735 26.375 8.525 28.255 ;
        RECT 96.540 13.245 97.555 14.080 ;
        RECT 63.980 8.230 65.740 9.725 ;
        RECT 156.660 1.440 157.100 1.880 ;
      LAYER met2 ;
        RECT 5.860 25.430 9.370 29.165 ;
        RECT 96.225 13.095 97.890 14.265 ;
        RECT 63.165 7.580 66.365 10.370 ;
        RECT 156.420 1.320 157.310 2.060 ;
      LAYER via2 ;
        RECT 6.735 26.375 8.525 28.255 ;
        RECT 96.540 13.245 97.555 14.080 ;
        RECT 63.980 8.230 65.740 9.725 ;
        RECT 156.660 1.440 157.100 1.880 ;
      LAYER met3 ;
        RECT 5.860 25.430 9.370 29.165 ;
        RECT 96.225 13.095 97.890 14.265 ;
        RECT 63.165 7.580 66.365 10.370 ;
        RECT 156.420 1.320 157.310 2.060 ;
      LAYER via3 ;
        RECT 6.735 26.375 8.525 28.255 ;
        RECT 96.540 13.245 97.555 14.080 ;
        RECT 63.980 8.230 65.740 9.725 ;
        RECT 156.660 1.440 157.100 1.880 ;
      LAYER met4 ;
        RECT 1.000 28.150 2.500 220.760 ;
        RECT 5.860 28.150 9.370 29.165 ;
        RECT 1.000 26.755 9.370 28.150 ;
        RECT 1.000 5.000 2.500 26.755 ;
        RECT 5.860 25.430 9.370 26.755 ;
        RECT 61.125 11.555 85.735 31.165 ;
        RECT 96.225 13.095 97.890 14.265 ;
        RECT 63.960 10.370 65.375 11.555 ;
        RECT 84.775 10.655 85.735 11.555 ;
        RECT 96.540 10.655 97.560 13.095 ;
        RECT 84.775 10.640 97.560 10.655 ;
        RECT 63.165 7.580 66.365 10.370 ;
        RECT 84.775 9.840 97.525 10.640 ;
        RECT 156.420 1.320 157.310 2.060 ;
        RECT 156.560 0.000 157.160 1.320 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 102.840 18.845 103.285 19.215 ;
        RECT 102.945 18.550 103.165 18.845 ;
        RECT 102.300 18.380 103.840 18.550 ;
      LAYER mcon ;
        RECT 102.955 18.925 103.150 19.150 ;
        RECT 102.380 18.380 103.760 18.550 ;
      LAYER met1 ;
        RECT 102.840 19.160 103.285 19.215 ;
        RECT 102.840 19.155 124.870 19.160 ;
        RECT 102.840 18.955 134.920 19.155 ;
        RECT 102.840 18.845 103.285 18.955 ;
        RECT 124.515 18.950 134.920 18.955 ;
        RECT 102.320 18.350 103.820 18.580 ;
        RECT 134.615 2.260 134.920 18.950 ;
        RECT 134.280 1.520 135.300 2.260 ;
      LAYER via ;
        RECT 134.490 1.650 135.090 2.110 ;
      LAYER met2 ;
        RECT 134.280 1.520 135.300 2.260 ;
      LAYER via2 ;
        RECT 134.490 1.650 135.090 2.110 ;
      LAYER met3 ;
        RECT 134.280 1.520 135.300 2.260 ;
      LAYER via3 ;
        RECT 134.490 1.650 135.090 2.110 ;
      LAYER met4 ;
        RECT 134.280 1.520 135.300 2.260 ;
        RECT 134.480 0.000 135.080 1.520 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER li1 ;
        RECT 88.600 22.300 89.260 22.700 ;
      LAYER mcon ;
        RECT 88.700 22.370 89.220 22.620 ;
      LAYER met1 ;
        RECT 88.595 22.300 89.265 22.705 ;
      LAYER via ;
        RECT 88.700 22.370 89.220 22.635 ;
      LAYER met2 ;
        RECT 88.595 22.300 89.265 22.705 ;
        RECT 88.735 20.240 88.945 22.300 ;
        RECT 88.735 20.055 88.950 20.240 ;
        RECT 88.740 15.155 88.950 20.055 ;
        RECT 88.740 14.805 112.890 15.155 ;
        RECT 88.740 14.800 88.950 14.805 ;
        RECT 112.540 2.310 112.890 14.805 ;
        RECT 112.210 1.435 113.215 2.310 ;
      LAYER via2 ;
        RECT 112.470 1.615 112.965 2.110 ;
      LAYER met3 ;
        RECT 112.210 1.435 113.215 2.310 ;
      LAYER via3 ;
        RECT 112.470 1.615 112.965 2.110 ;
      LAYER met4 ;
        RECT 112.210 1.435 113.215 2.310 ;
        RECT 112.395 0.905 113.005 1.435 ;
        RECT 112.400 0.000 113.000 0.905 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 89.480 22.175 91.520 22.345 ;
        RECT 89.500 21.440 91.500 22.175 ;
        RECT 93.630 21.800 95.170 21.970 ;
        RECT 89.510 15.830 91.500 21.440 ;
        RECT 93.645 20.840 95.150 21.800 ;
        RECT 102.295 21.790 103.135 21.960 ;
        RECT 104.745 21.850 106.285 22.020 ;
        RECT 102.630 21.135 102.800 21.790 ;
        RECT 93.700 15.830 95.060 20.840 ;
        RECT 102.560 20.785 102.905 21.135 ;
        RECT 104.765 21.020 106.265 21.850 ;
        RECT 98.520 17.895 100.060 18.065 ;
        RECT 98.540 17.070 100.040 17.895 ;
        RECT 98.550 15.830 100.035 17.070 ;
        RECT 104.770 15.830 106.260 21.020 ;
        RECT 88.710 13.075 90.500 14.225 ;
        RECT 88.915 11.790 90.330 13.075 ;
        RECT 88.915 10.375 107.255 11.790 ;
        RECT 105.840 9.615 107.255 10.375 ;
        RECT 105.335 8.205 107.495 9.615 ;
      LAYER mcon ;
        RECT 89.560 22.175 91.440 22.345 ;
        RECT 93.710 21.800 95.090 21.970 ;
        RECT 102.375 21.790 103.055 21.960 ;
        RECT 104.825 21.850 106.205 22.020 ;
        RECT 102.640 20.860 102.815 21.035 ;
        RECT 89.805 16.020 91.170 16.425 ;
        RECT 98.600 17.895 99.980 18.065 ;
        RECT 94.000 16.070 94.770 16.460 ;
        RECT 98.705 16.020 99.855 16.440 ;
        RECT 105.195 16.035 105.895 16.490 ;
        RECT 89.060 13.270 90.165 14.045 ;
        RECT 105.420 8.285 107.405 9.535 ;
      LAYER met1 ;
        RECT 89.500 22.145 91.500 22.375 ;
        RECT 93.650 21.770 95.150 22.000 ;
        RECT 102.315 21.760 103.115 21.990 ;
        RECT 104.765 21.820 106.265 22.050 ;
        RECT 102.560 20.785 102.905 21.135 ;
        RECT 102.615 20.600 102.855 20.785 ;
        RECT 101.350 20.360 102.855 20.600 ;
        RECT 98.540 17.865 100.040 18.095 ;
        RECT 51.520 16.610 53.095 16.950 ;
        RECT 101.350 16.610 101.590 20.360 ;
        RECT 51.520 16.600 54.295 16.610 ;
        RECT 88.710 16.600 106.270 16.610 ;
        RECT 51.520 15.830 106.270 16.600 ;
        RECT 51.520 15.815 90.500 15.830 ;
        RECT 51.520 15.550 53.095 15.815 ;
        RECT 88.710 13.075 90.500 15.815 ;
        RECT 105.360 8.255 107.465 9.565 ;
      LAYER via ;
        RECT 51.840 15.840 52.760 16.670 ;
        RECT 89.060 13.270 90.165 14.045 ;
      LAYER met2 ;
        RECT 51.520 15.550 53.095 16.950 ;
        RECT 88.710 13.075 90.500 14.225 ;
      LAYER via2 ;
        RECT 51.840 15.840 52.760 16.670 ;
        RECT 89.060 13.270 90.165 14.045 ;
      LAYER met3 ;
        RECT 51.520 15.550 53.095 16.950 ;
        RECT 60.730 13.785 87.590 31.560 ;
        RECT 88.710 13.785 90.500 14.225 ;
        RECT 60.730 13.370 90.500 13.785 ;
        RECT 60.730 11.160 87.590 13.370 ;
        RECT 88.710 13.075 90.500 13.370 ;
      LAYER via3 ;
        RECT 51.840 15.840 52.760 16.670 ;
        RECT 87.170 11.300 87.490 31.420 ;
      LAYER met4 ;
        RECT 49.000 16.610 50.500 220.760 ;
        RECT 51.520 16.610 53.095 16.950 ;
        RECT 49.000 15.815 53.095 16.610 ;
        RECT 49.000 5.000 50.500 15.815 ;
        RECT 51.520 15.550 53.095 15.815 ;
        RECT 87.090 11.220 87.570 31.500 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 103.705 24.495 104.035 24.560 ;
        RECT 104.330 24.495 104.540 24.500 ;
        RECT 103.705 24.325 104.540 24.495 ;
        RECT 88.850 24.060 92.130 24.230 ;
        RECT 103.705 24.220 104.035 24.325 ;
        RECT 89.565 23.465 91.445 24.060 ;
        RECT 92.410 23.650 92.745 23.925 ;
        RECT 92.470 23.465 92.685 23.650 ;
        RECT 89.565 23.280 92.685 23.465 ;
        RECT 89.565 22.815 91.445 23.280 ;
        RECT 104.330 22.930 104.540 24.325 ;
        RECT 89.480 22.645 91.520 22.815 ;
        RECT 103.660 22.760 104.540 22.930 ;
        RECT 101.805 21.940 102.120 22.275 ;
        RECT 97.620 21.570 100.900 21.740 ;
        RECT 98.520 21.290 99.900 21.570 ;
        RECT 98.520 21.115 100.725 21.290 ;
        RECT 98.520 20.915 99.900 21.115 ;
        RECT 98.470 20.745 100.010 20.915 ;
        RECT 100.555 20.750 100.725 21.115 ;
        RECT 100.555 20.560 100.730 20.750 ;
        RECT 98.470 20.275 100.010 20.445 ;
        RECT 98.490 19.470 99.990 20.275 ;
        RECT 100.560 20.190 100.730 20.560 ;
        RECT 101.875 20.190 102.055 21.940 ;
        RECT 103.660 20.190 103.890 22.760 ;
        RECT 104.330 22.390 104.540 22.760 ;
        RECT 104.190 21.990 104.560 22.390 ;
        RECT 100.560 20.020 103.890 20.190 ;
        RECT 98.635 19.105 99.850 19.470 ;
        RECT 98.635 19.095 101.255 19.105 ;
        RECT 98.635 18.925 101.260 19.095 ;
        RECT 98.635 18.535 99.850 18.925 ;
        RECT 98.520 18.365 100.060 18.535 ;
        RECT 101.055 17.440 101.260 18.925 ;
        RECT 101.875 18.425 102.065 20.020 ;
        RECT 102.275 20.015 103.695 20.020 ;
        RECT 101.845 18.045 102.120 18.425 ;
        RECT 102.300 17.910 103.840 18.080 ;
        RECT 102.315 17.440 103.825 17.910 ;
        RECT 101.055 17.255 103.825 17.440 ;
        RECT 102.315 17.070 103.825 17.255 ;
      LAYER mcon ;
        RECT 88.930 24.060 92.050 24.230 ;
        RECT 89.560 22.645 91.440 22.815 ;
        RECT 97.700 21.570 100.820 21.740 ;
        RECT 98.550 20.745 99.930 20.915 ;
        RECT 98.550 20.275 99.930 20.445 ;
        RECT 98.600 18.365 99.980 18.535 ;
        RECT 102.380 17.910 103.760 18.080 ;
      LAYER met1 ;
        RECT 88.870 24.030 92.110 24.260 ;
        RECT 89.500 22.615 91.500 22.845 ;
        RECT 97.640 21.540 100.880 21.770 ;
        RECT 98.490 20.715 99.990 20.945 ;
        RECT 98.490 20.245 99.990 20.475 ;
        RECT 98.540 18.335 100.040 18.565 ;
        RECT 102.320 17.880 103.820 18.110 ;
  END
END tt_um_analog_example
END LIBRARY

