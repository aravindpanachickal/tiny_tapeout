magic
tech sky130B
magscale 1 2
timestamp 1713363624
<< poly >>
rect 17720 4460 17852 4540
<< locali >>
rect 17720 4524 17852 4540
rect 17720 4474 17740 4524
rect 17844 4474 17852 4524
rect 17720 4460 17852 4474
<< viali >>
rect 17740 4474 17844 4524
<< metal1 >>
rect 1172 5651 1874 5833
rect 1172 5275 1347 5651
rect 1705 5634 1874 5651
rect 17659 5634 17763 5635
rect 1705 5354 17939 5634
rect 1705 5275 1874 5354
rect 17659 5352 17763 5354
rect 1172 5086 1874 5275
rect 21538 4680 31404 4710
rect 17719 4527 17853 4541
rect 17719 4474 17740 4527
rect 17844 4474 17853 4527
rect 17719 4460 17853 4474
rect 21414 3831 24974 3832
rect 21414 3791 26984 3831
rect 24903 3790 26984 3791
rect 10304 3334 10619 3390
rect 10304 3168 10368 3334
rect 10552 3322 10619 3334
rect 10552 3320 10859 3322
rect 10552 3168 17815 3320
rect 10304 3163 17815 3168
rect 10304 3110 10619 3163
rect 26923 452 26984 3790
rect 26856 422 27060 452
rect 26856 330 26898 422
rect 27018 330 27060 422
rect 31346 412 31404 4680
rect 26856 304 27060 330
rect 31284 376 31462 412
rect 31284 288 31332 376
rect 31420 288 31462 376
rect 31284 264 31462 288
<< via1 >>
rect 1347 5275 1705 5651
rect 17740 4524 17844 4527
rect 17740 4474 17844 4524
rect 10368 3168 10552 3334
rect 26898 330 27018 422
rect 31332 288 31420 376
<< metal2 >>
rect 1172 5651 1874 5833
rect 1172 5275 1347 5651
rect 1705 5275 1874 5651
rect 1172 5086 1874 5275
rect 17719 4527 17853 4541
rect 17719 4474 17740 4527
rect 17844 4474 17853 4527
rect 17719 4460 17853 4474
rect 17747 4048 17789 4460
rect 17747 4011 17790 4048
rect 10304 3334 10619 3390
rect 10304 3168 10368 3334
rect 10552 3168 10619 3334
rect 10304 3110 10619 3168
rect 17748 3031 17790 4011
rect 17748 2961 22578 3031
rect 17748 2960 17790 2961
rect 22508 462 22578 2961
rect 22442 422 22643 462
rect 22442 323 22494 422
rect 22593 323 22643 422
rect 22442 287 22643 323
rect 26856 422 27060 452
rect 26856 330 26898 422
rect 27018 330 27060 422
rect 26856 304 27060 330
rect 31284 376 31462 412
rect 31284 288 31332 376
rect 31420 288 31462 376
rect 31284 264 31462 288
<< via2 >>
rect 1347 5275 1705 5651
rect 10368 3168 10552 3334
rect 22494 323 22593 422
rect 26898 330 27018 422
rect 31332 288 31420 376
<< metal3 >>
rect 1172 5651 1874 5833
rect 1172 5275 1347 5651
rect 1705 5275 1874 5651
rect 1172 5086 1874 5275
rect 10304 3334 10619 3390
rect 10304 3168 10368 3334
rect 10552 3168 10619 3334
rect 10304 3110 10619 3168
rect 22442 422 22643 462
rect 22442 323 22494 422
rect 22593 323 22643 422
rect 22442 287 22643 323
rect 26856 422 27060 452
rect 26856 330 26898 422
rect 27018 330 27060 422
rect 26856 304 27060 330
rect 31284 376 31462 412
rect 31284 288 31332 376
rect 31420 288 31462 376
rect 31284 264 31462 288
<< via3 >>
rect 1347 5275 1705 5651
rect 10368 3168 10552 3334
rect 22494 323 22593 422
rect 26898 330 27018 422
rect 31332 288 31420 376
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 5630 500 44152
rect 1172 5651 1874 5833
rect 1172 5630 1347 5651
rect 200 5351 1347 5630
rect 200 1000 500 5351
rect 1172 5275 1347 5351
rect 1705 5275 1874 5651
rect 1172 5086 1874 5275
rect 9800 3322 10100 44152
rect 10304 3334 10619 3390
rect 10304 3322 10368 3334
rect 9800 3168 10368 3322
rect 10552 3168 10619 3334
rect 9800 3163 10619 3168
rect 9800 1000 10100 3163
rect 10304 3110 10619 3163
rect 22442 422 22643 462
rect 22442 323 22494 422
rect 22593 323 22643 422
rect 22442 287 22643 323
rect 26856 422 27060 452
rect 26856 330 26898 422
rect 27018 330 27060 422
rect 26856 304 27060 330
rect 31284 376 31462 412
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22479 181 22601 287
rect 22480 0 22600 181
rect 26896 0 27016 304
rect 31284 288 31332 376
rect 31420 288 31462 376
rect 31284 264 31462 288
rect 31312 0 31432 264
use leakylayout  leakylayout_0 ~/Desktop/workbench/SNN/simulation/leaky.sch
timestamp 1713357858
transform 1 0 18302 0 1 2824
box -6156 -1308 3342 3488
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
