magic
tech sky130A
timestamp 1713438817
<< error_p >>
rect -56 -91 56 91
<< nwell >>
rect -56 -91 56 91
<< pmos >>
rect -9 -60 9 60
<< pdiff >>
rect -38 54 -9 60
rect -38 -54 -32 54
rect -15 -54 -9 54
rect -38 -60 -9 -54
rect 9 54 38 60
rect 9 -54 15 54
rect 32 -54 38 54
rect 9 -60 38 -54
<< pdiffc >>
rect -32 -54 -15 54
rect 15 -54 32 54
<< poly >>
rect -9 60 9 73
rect -9 -73 9 -60
<< locali >>
rect -32 54 -15 62
rect -32 -62 -15 -54
rect 15 54 32 62
rect 15 -62 32 -54
<< viali >>
rect -32 -54 -15 54
rect 15 -54 32 54
<< metal1 >>
rect -35 54 -12 60
rect -35 -54 -32 54
rect -15 -54 -12 54
rect -35 -60 -12 -54
rect 12 54 35 60
rect 12 -54 15 54
rect 32 -54 35 54
rect 12 -60 35 -54
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.2 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
