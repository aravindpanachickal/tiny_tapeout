VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO leakylayout
  CLASS BLOCK ;
  FOREIGN leakylayout ;
  ORIGIN 30.780 6.540 ;
  SIZE 47.490 BY 23.980 ;
  OBS
      LAYER nwell ;
        RECT -2.950 9.650 12.780 12.600 ;
        RECT 0.620 9.465 1.495 9.650 ;
        RECT 5.240 9.445 12.780 9.650 ;
        RECT 5.240 7.915 12.765 9.445 ;
        RECT 5.240 7.150 12.760 7.915 ;
        RECT 5.240 7.140 10.010 7.150 ;
      LAYER li1 ;
        RECT -2.645 10.580 0.605 14.050 ;
        RECT 1.580 10.585 4.830 14.050 ;
        RECT -2.660 10.410 0.620 10.580 ;
        RECT 1.570 10.415 4.850 10.585 ;
        RECT 6.040 10.580 9.290 14.050 ;
        RECT -2.660 9.940 0.620 10.110 ;
        RECT 1.570 9.945 4.850 10.115 ;
        RECT 5.425 10.040 5.760 10.465 ;
        RECT 6.020 10.410 9.300 10.580 ;
        RECT 10.660 10.575 11.860 14.050 ;
        RECT 10.640 10.405 11.880 10.575 ;
        RECT 12.195 10.375 12.525 10.440 ;
        RECT 12.820 10.375 13.030 10.380 ;
        RECT 12.195 10.205 13.030 10.375 ;
        RECT -1.945 9.345 -0.065 9.940 ;
        RECT 0.900 9.530 1.235 9.805 ;
        RECT 0.960 9.345 1.175 9.530 ;
        RECT -1.945 9.160 1.175 9.345 ;
        RECT 2.745 9.340 3.125 9.945 ;
        RECT 2.745 9.325 4.945 9.340 ;
        RECT -1.945 8.695 -0.065 9.160 ;
        RECT 2.745 9.090 4.955 9.325 ;
        RECT -2.555 8.455 -2.255 8.575 ;
        RECT -2.030 8.525 0.010 8.695 ;
        RECT -2.910 8.275 -2.255 8.455 ;
        RECT 4.740 8.320 4.955 9.090 ;
        RECT -2.555 8.180 -2.255 8.275 ;
        RECT -2.030 8.055 0.010 8.225 ;
        RECT -2.010 7.320 -0.010 8.055 ;
        RECT 1.440 7.745 1.900 8.225 ;
        RECT 2.120 8.150 4.960 8.320 ;
        RECT 2.120 7.680 3.660 7.850 ;
        RECT -2.000 1.710 -0.010 7.320 ;
        RECT 2.135 6.720 3.640 7.680 ;
        RECT 4.740 6.995 4.955 8.150 ;
        RECT 5.525 7.955 5.695 10.040 ;
        RECT 6.020 9.940 9.300 10.110 ;
        RECT 6.385 9.660 9.180 9.940 ;
        RECT 10.640 9.935 11.880 10.105 ;
        RECT 12.195 10.100 12.525 10.205 ;
        RECT 11.135 9.740 11.305 9.935 ;
        RECT 6.385 9.490 10.255 9.660 ;
        RECT 11.130 9.535 11.305 9.740 ;
        RECT 6.385 9.300 9.180 9.490 ;
        RECT 6.130 8.090 9.370 9.300 ;
        RECT 10.085 8.905 10.255 9.490 ;
        RECT 11.065 9.195 11.390 9.535 ;
        RECT 10.085 8.900 11.595 8.905 ;
        RECT 10.085 8.735 11.605 8.900 ;
        RECT 12.820 8.810 13.030 10.205 ;
        RECT 10.805 8.310 11.605 8.735 ;
        RECT 12.150 8.640 13.030 8.810 ;
        RECT 5.430 7.560 5.805 7.955 ;
        RECT 6.110 7.920 9.390 8.090 ;
        RECT 10.295 7.820 10.610 8.155 ;
        RECT 10.785 8.140 11.625 8.310 ;
        RECT 5.540 6.995 5.710 7.560 ;
        RECT 6.110 7.450 9.390 7.620 ;
        RECT 7.010 7.170 8.390 7.450 ;
        RECT 7.010 6.995 9.215 7.170 ;
        RECT 4.740 6.815 5.715 6.995 ;
        RECT 4.755 6.810 5.715 6.815 ;
        RECT 2.190 1.710 3.550 6.720 ;
        RECT 5.540 6.540 5.710 6.810 ;
        RECT 7.010 6.730 8.390 6.995 ;
        RECT 5.535 6.500 5.710 6.540 ;
        RECT 6.335 6.500 6.640 6.580 ;
        RECT 6.960 6.560 8.500 6.730 ;
        RECT 9.045 6.630 9.215 6.995 ;
        RECT 5.535 6.330 6.640 6.500 ;
        RECT 9.045 6.440 9.220 6.630 ;
        RECT 5.535 4.185 5.710 6.330 ;
        RECT 6.335 6.225 6.640 6.330 ;
        RECT 6.960 6.090 8.500 6.260 ;
        RECT 6.980 5.285 8.480 6.090 ;
        RECT 9.050 6.070 9.220 6.440 ;
        RECT 10.365 6.070 10.545 7.820 ;
        RECT 10.785 7.670 11.625 7.840 ;
        RECT 11.120 7.015 11.290 7.670 ;
        RECT 11.050 6.665 11.395 7.015 ;
        RECT 12.150 6.070 12.380 8.640 ;
        RECT 12.820 8.270 13.030 8.640 ;
        RECT 13.695 8.605 14.140 8.975 ;
        RECT 13.800 8.370 14.010 8.605 ;
        RECT 12.680 7.870 13.050 8.270 ;
        RECT 13.235 8.200 14.775 8.370 ;
        RECT 13.235 7.730 14.775 7.900 ;
        RECT 13.255 6.900 14.755 7.730 ;
        RECT 9.050 5.900 12.380 6.070 ;
        RECT 7.125 4.985 8.340 5.285 ;
        RECT 7.125 4.975 9.745 4.985 ;
        RECT 7.125 4.805 9.750 4.975 ;
        RECT 7.125 4.415 8.340 4.805 ;
        RECT 6.455 4.185 6.795 4.280 ;
        RECT 7.010 4.245 8.550 4.415 ;
        RECT 5.535 4.010 6.795 4.185 ;
        RECT 5.535 0.145 5.750 4.010 ;
        RECT 6.455 3.930 6.795 4.010 ;
        RECT 7.010 3.775 8.550 3.945 ;
        RECT 7.030 2.950 8.530 3.775 ;
        RECT 9.545 3.320 9.750 4.805 ;
        RECT 10.365 4.305 10.555 5.900 ;
        RECT 10.765 5.895 12.185 5.900 ;
        RECT 11.330 4.725 11.775 5.095 ;
        RECT 11.435 4.430 11.655 4.725 ;
        RECT 10.335 3.925 10.610 4.305 ;
        RECT 10.790 4.260 12.330 4.430 ;
        RECT 10.790 3.790 12.330 3.960 ;
        RECT 10.805 3.320 12.315 3.790 ;
        RECT 9.545 3.135 12.315 3.320 ;
        RECT 10.805 2.950 12.315 3.135 ;
        RECT 7.040 1.710 8.525 2.950 ;
        RECT 13.260 1.710 14.750 6.900 ;
        RECT -2.800 -1.045 -1.010 0.105 ;
        RECT 4.715 -1.025 6.380 0.145 ;
        RECT -2.595 -2.330 -1.180 -1.045 ;
        RECT -2.595 -3.745 15.745 -2.330 ;
        RECT -28.345 -4.505 -25.145 -3.750 ;
        RECT 14.330 -4.505 15.745 -3.745 ;
        RECT -28.345 -5.915 -21.615 -4.505 ;
        RECT 13.825 -5.915 15.985 -4.505 ;
        RECT -28.345 -6.540 -25.145 -5.915 ;
      LAYER mcon ;
        RECT -1.445 12.970 -0.610 13.725 ;
        RECT 2.830 12.960 3.665 13.715 ;
        RECT 7.220 12.955 8.055 13.710 ;
        RECT -2.580 10.410 0.540 10.580 ;
        RECT 1.650 10.415 4.770 10.585 ;
        RECT 10.865 12.935 11.700 13.690 ;
        RECT -2.580 9.940 0.540 10.110 ;
        RECT 1.650 9.945 4.770 10.115 ;
        RECT 6.100 10.410 9.220 10.580 ;
        RECT 10.720 10.405 11.800 10.575 ;
        RECT -1.950 8.525 -0.070 8.695 ;
        RECT -1.950 8.055 -0.070 8.225 ;
        RECT 1.500 7.830 1.850 8.160 ;
        RECT 2.200 8.150 3.580 8.320 ;
        RECT 2.200 7.680 3.580 7.850 ;
        RECT 6.100 9.940 9.220 10.110 ;
        RECT 10.720 9.935 11.800 10.105 ;
        RECT 11.125 9.250 11.325 9.460 ;
        RECT 6.190 7.920 9.310 8.090 ;
        RECT 10.865 8.140 11.545 8.310 ;
        RECT 6.190 7.450 9.310 7.620 ;
        RECT -1.705 1.900 -0.340 2.305 ;
        RECT 2.490 1.950 3.260 2.340 ;
        RECT 7.040 6.560 8.420 6.730 ;
        RECT 7.040 6.090 8.420 6.260 ;
        RECT 10.865 7.670 11.545 7.840 ;
        RECT 11.130 6.740 11.305 6.915 ;
        RECT 13.825 8.695 14.035 8.880 ;
        RECT 13.315 8.200 14.695 8.370 ;
        RECT 13.315 7.730 14.695 7.900 ;
        RECT 7.090 4.245 8.470 4.415 ;
        RECT 7.090 3.775 8.470 3.945 ;
        RECT 11.445 4.805 11.640 5.030 ;
        RECT 10.870 4.260 12.250 4.430 ;
        RECT 10.870 3.790 12.250 3.960 ;
        RECT 7.195 1.900 8.345 2.320 ;
        RECT 13.685 1.915 14.385 2.370 ;
        RECT -2.450 -0.850 -1.345 -0.075 ;
        RECT 5.030 -0.875 6.045 -0.040 ;
        RECT -27.530 -5.890 -25.770 -4.395 ;
        RECT -23.685 -5.835 -21.700 -4.585 ;
        RECT 13.910 -5.835 15.895 -4.585 ;
      LAYER met1 ;
        RECT -2.950 12.650 12.735 14.050 ;
        RECT 1.575 11.920 15.425 12.105 ;
        RECT 1.580 11.065 1.745 11.920 ;
        RECT 1.585 10.615 1.745 11.065 ;
        RECT -2.640 10.380 0.600 10.610 ;
        RECT 1.585 10.385 4.830 10.615 ;
        RECT 1.585 10.145 1.745 10.385 ;
        RECT 6.040 10.380 9.280 10.610 ;
        RECT 10.660 10.375 11.860 10.605 ;
        RECT -2.640 9.910 0.600 10.140 ;
        RECT 1.585 9.915 4.830 10.145 ;
        RECT -2.010 8.495 -0.010 8.725 ;
        RECT 1.585 8.310 1.745 9.915 ;
        RECT 6.040 9.910 9.280 10.140 ;
        RECT 10.660 9.905 11.860 10.135 ;
        RECT 11.065 9.430 11.390 9.535 ;
        RECT 15.255 9.430 15.425 11.920 ;
        RECT 11.065 9.290 16.710 9.430 ;
        RECT 11.065 9.285 15.425 9.290 ;
        RECT 15.775 9.285 16.710 9.290 ;
        RECT 11.065 9.195 11.390 9.285 ;
        RECT 13.850 8.975 13.990 9.285 ;
        RECT 13.695 8.605 14.140 8.975 ;
        RECT -2.010 8.025 -0.010 8.255 ;
        RECT 1.360 7.645 1.975 8.310 ;
        RECT 2.140 8.120 3.640 8.350 ;
        RECT 6.130 7.890 9.370 8.120 ;
        RECT 10.805 8.110 11.605 8.340 ;
        RECT 13.255 8.170 14.755 8.400 ;
        RECT 2.140 7.650 3.640 7.880 ;
        RECT 1.585 7.640 1.800 7.645 ;
        RECT 6.130 7.420 9.370 7.650 ;
        RECT 10.805 7.640 11.605 7.870 ;
        RECT 13.255 7.700 14.755 7.930 ;
        RECT 6.980 6.530 8.480 6.760 ;
        RECT 11.050 6.665 11.395 7.015 ;
        RECT 11.105 6.480 11.345 6.665 ;
        RECT 6.980 6.060 8.480 6.290 ;
        RECT 9.840 6.240 11.345 6.480 ;
        RECT 7.030 4.215 8.530 4.445 ;
        RECT 7.030 3.745 8.530 3.975 ;
        RECT 9.840 2.490 10.080 6.240 ;
        RECT 11.330 5.040 11.775 5.095 ;
        RECT 11.330 4.835 15.970 5.040 ;
        RECT 11.330 4.725 11.775 4.835 ;
        RECT 10.810 4.230 12.310 4.460 ;
        RECT 10.810 3.760 12.310 3.990 ;
        RECT -2.800 1.710 14.760 2.490 ;
        RECT -2.800 -1.045 -1.010 1.710 ;
        RECT 4.715 -1.025 6.380 0.145 ;
        RECT -28.345 -6.540 -25.145 -3.750 ;
        RECT -23.745 -5.865 -21.640 -4.555 ;
        RECT 13.850 -5.865 15.955 -4.555 ;
      LAYER via ;
        RECT -2.450 -0.850 -1.345 -0.075 ;
        RECT 5.030 -0.875 6.045 -0.040 ;
        RECT -27.530 -5.890 -25.770 -4.395 ;
      LAYER met2 ;
        RECT -2.800 -1.045 -1.010 0.105 ;
        RECT 4.715 -1.025 6.380 0.145 ;
        RECT -28.345 -6.540 -25.145 -3.750 ;
      LAYER via2 ;
        RECT -2.450 -0.850 -1.345 -0.075 ;
        RECT 5.030 -0.875 6.045 -0.040 ;
        RECT -27.530 -5.890 -25.770 -4.395 ;
      LAYER met3 ;
        RECT -30.780 -0.335 -3.920 17.440 ;
        RECT -2.710 -0.335 -1.010 0.105 ;
        RECT -30.780 -0.750 -1.010 -0.335 ;
        RECT -30.780 -2.960 -3.920 -0.750 ;
        RECT -2.710 -1.045 -1.010 -0.750 ;
        RECT 4.715 -1.025 6.380 0.145 ;
        RECT -28.345 -6.540 -25.145 -3.750 ;
      LAYER via3 ;
        RECT -4.340 -2.820 -4.020 17.300 ;
        RECT 5.030 -0.875 6.045 -0.040 ;
        RECT -27.530 -5.890 -25.770 -4.395 ;
      LAYER met4 ;
        RECT -30.385 -2.565 -5.775 17.045 ;
        RECT -27.550 -3.750 -26.135 -2.565 ;
        RECT -6.735 -3.465 -5.775 -2.565 ;
        RECT -4.420 -2.900 -3.940 17.380 ;
        RECT 4.715 -1.025 6.380 0.145 ;
        RECT 5.030 -3.465 6.050 -1.025 ;
        RECT -6.735 -3.480 6.050 -3.465 ;
        RECT -28.345 -6.540 -25.145 -3.750 ;
        RECT -6.735 -4.280 6.015 -3.480 ;
  END
END leakylayout
END LIBRARY

