VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_lif
  CLASS BLOCK ;
  FOREIGN tt_um_lif ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.976400 ;
    ANTENNADIFFAREA 28.198374 ;
    PORT
      LAYER nwell ;
        RECT 85.040 23.650 100.770 26.600 ;
        RECT 88.610 23.465 89.485 23.650 ;
        RECT 93.230 23.445 100.770 23.650 ;
        RECT 93.230 21.915 100.755 23.445 ;
        RECT 93.230 21.150 100.750 21.915 ;
        RECT 93.230 21.140 98.000 21.150 ;
      LAYER li1 ;
        RECT 85.345 24.580 88.595 28.050 ;
        RECT 89.570 24.585 92.820 28.050 ;
        RECT 85.330 24.410 88.610 24.580 ;
        RECT 89.560 24.415 92.840 24.585 ;
        RECT 94.030 24.580 97.280 28.050 ;
        RECT 89.560 23.945 92.840 24.115 ;
        RECT 93.415 24.040 93.750 24.465 ;
        RECT 94.010 24.410 97.290 24.580 ;
        RECT 98.650 24.575 99.850 28.050 ;
        RECT 98.630 24.405 99.870 24.575 ;
        RECT 90.735 23.340 91.115 23.945 ;
        RECT 90.735 23.325 92.935 23.340 ;
        RECT 90.735 23.090 92.945 23.325 ;
        RECT 92.730 22.320 92.945 23.090 ;
        RECT 89.430 21.745 89.890 22.225 ;
        RECT 90.110 22.150 92.950 22.320 ;
        RECT 92.730 20.995 92.945 22.150 ;
        RECT 93.515 21.955 93.685 24.040 ;
        RECT 94.010 23.940 97.290 24.110 ;
        RECT 94.375 23.660 97.170 23.940 ;
        RECT 98.630 23.935 99.870 24.105 ;
        RECT 99.125 23.740 99.295 23.935 ;
        RECT 94.375 23.490 98.245 23.660 ;
        RECT 99.120 23.535 99.295 23.740 ;
        RECT 94.375 23.300 97.170 23.490 ;
        RECT 94.120 22.090 97.360 23.300 ;
        RECT 98.075 22.905 98.245 23.490 ;
        RECT 99.055 23.195 99.380 23.535 ;
        RECT 98.075 22.900 99.585 22.905 ;
        RECT 98.075 22.735 99.595 22.900 ;
        RECT 98.795 22.310 99.595 22.735 ;
        RECT 101.685 22.605 102.130 22.975 ;
        RECT 101.790 22.370 102.000 22.605 ;
        RECT 98.775 22.140 99.615 22.310 ;
        RECT 101.225 22.200 102.765 22.370 ;
        RECT 93.420 21.560 93.795 21.955 ;
        RECT 94.100 21.920 97.380 22.090 ;
        RECT 93.530 20.995 93.700 21.560 ;
        RECT 92.730 20.815 93.705 20.995 ;
        RECT 92.745 20.810 93.705 20.815 ;
        RECT 93.530 20.540 93.700 20.810 ;
        RECT 93.525 20.500 93.700 20.540 ;
        RECT 94.325 20.500 94.630 20.580 ;
        RECT 93.525 20.330 94.630 20.500 ;
        RECT 93.525 18.185 93.700 20.330 ;
        RECT 94.325 20.225 94.630 20.330 ;
        RECT 94.445 18.185 94.785 18.280 ;
        RECT 93.525 18.010 94.785 18.185 ;
        RECT 93.525 14.145 93.740 18.010 ;
        RECT 94.445 17.930 94.785 18.010 ;
        RECT 92.705 12.975 94.370 14.145 ;
        RECT 59.645 9.495 62.845 10.250 ;
        RECT 59.645 8.085 66.375 9.495 ;
        RECT 59.645 7.460 62.845 8.085 ;
      LAYER mcon ;
        RECT 86.545 26.970 87.380 27.725 ;
        RECT 90.820 26.960 91.655 27.715 ;
        RECT 95.210 26.955 96.045 27.710 ;
        RECT 85.410 24.410 88.530 24.580 ;
        RECT 89.640 24.415 92.760 24.585 ;
        RECT 98.855 26.935 99.690 27.690 ;
        RECT 89.640 23.945 92.760 24.115 ;
        RECT 94.090 24.410 97.210 24.580 ;
        RECT 98.710 24.405 99.790 24.575 ;
        RECT 89.490 21.830 89.840 22.160 ;
        RECT 90.190 22.150 91.570 22.320 ;
        RECT 94.090 23.940 97.210 24.110 ;
        RECT 98.710 23.935 99.790 24.105 ;
        RECT 99.115 23.250 99.315 23.460 ;
        RECT 101.815 22.695 102.025 22.880 ;
        RECT 98.855 22.140 99.535 22.310 ;
        RECT 101.305 22.200 102.685 22.370 ;
        RECT 94.180 21.920 97.300 22.090 ;
        RECT 93.020 13.125 94.035 13.960 ;
        RECT 60.460 8.110 62.220 9.605 ;
        RECT 64.305 8.165 66.290 9.415 ;
      LAYER met1 ;
        RECT 4.210 28.050 7.175 28.775 ;
        RECT 4.210 26.650 100.725 28.050 ;
        RECT 4.210 26.225 7.175 26.650 ;
        RECT 89.565 25.920 103.415 26.105 ;
        RECT 89.570 25.065 89.735 25.920 ;
        RECT 89.575 24.615 89.735 25.065 ;
        RECT 85.350 24.380 88.590 24.610 ;
        RECT 89.575 24.385 92.820 24.615 ;
        RECT 89.575 24.145 89.735 24.385 ;
        RECT 94.030 24.380 97.270 24.610 ;
        RECT 98.650 24.375 99.850 24.605 ;
        RECT 89.575 23.915 92.820 24.145 ;
        RECT 89.575 22.310 89.735 23.915 ;
        RECT 94.030 23.910 97.270 24.140 ;
        RECT 98.650 23.905 99.850 24.135 ;
        RECT 99.055 23.430 99.380 23.535 ;
        RECT 103.245 23.430 103.415 25.920 ;
        RECT 99.055 23.290 156.920 23.430 ;
        RECT 99.055 23.285 103.415 23.290 ;
        RECT 103.765 23.285 156.920 23.290 ;
        RECT 99.055 23.195 99.380 23.285 ;
        RECT 101.840 22.975 101.980 23.285 ;
        RECT 101.685 22.605 102.130 22.975 ;
        RECT 89.350 21.645 89.965 22.310 ;
        RECT 90.130 22.120 91.630 22.350 ;
        RECT 94.120 21.890 97.360 22.120 ;
        RECT 98.795 22.110 99.595 22.340 ;
        RECT 101.245 22.170 102.745 22.400 ;
        RECT 89.575 21.640 89.790 21.645 ;
        RECT 92.705 12.975 94.370 14.145 ;
        RECT 59.645 7.460 62.845 10.250 ;
        RECT 64.245 8.135 66.350 9.445 ;
        RECT 156.775 2.280 156.915 23.285 ;
        RECT 156.490 1.620 157.260 2.280 ;
      LAYER via ;
        RECT 4.885 26.720 6.560 28.120 ;
        RECT 93.020 13.125 94.035 13.960 ;
        RECT 60.460 8.110 62.220 9.605 ;
        RECT 156.650 1.780 157.120 2.140 ;
      LAYER met2 ;
        RECT 4.210 26.225 7.175 28.775 ;
        RECT 92.705 12.975 94.370 14.145 ;
        RECT 59.645 7.460 62.845 10.250 ;
        RECT 156.490 1.620 157.260 2.280 ;
      LAYER via2 ;
        RECT 4.885 26.720 6.560 28.120 ;
        RECT 93.020 13.125 94.035 13.960 ;
        RECT 60.460 8.110 62.220 9.605 ;
        RECT 156.650 1.780 157.120 2.140 ;
      LAYER met3 ;
        RECT 4.210 26.225 7.175 28.775 ;
        RECT 92.705 12.975 94.370 14.145 ;
        RECT 59.645 7.460 62.845 10.250 ;
        RECT 156.490 1.620 157.260 2.280 ;
      LAYER via3 ;
        RECT 4.885 26.720 6.560 28.120 ;
        RECT 93.020 13.125 94.035 13.960 ;
        RECT 60.460 8.110 62.220 9.605 ;
        RECT 156.650 1.780 157.120 2.140 ;
      LAYER met4 ;
        RECT 1.000 28.040 2.500 220.760 ;
        RECT 4.210 28.040 7.175 28.775 ;
        RECT 1.000 26.655 7.175 28.040 ;
        RECT 1.000 5.000 2.500 26.655 ;
        RECT 4.210 26.225 7.175 26.655 ;
        RECT 57.605 11.435 82.215 31.045 ;
        RECT 92.705 12.975 94.370 14.145 ;
        RECT 60.440 10.250 61.855 11.435 ;
        RECT 81.255 10.535 82.215 11.435 ;
        RECT 93.020 10.535 94.040 12.975 ;
        RECT 81.255 10.520 94.040 10.535 ;
        RECT 59.645 7.460 62.845 10.250 ;
        RECT 81.255 9.720 94.005 10.520 ;
        RECT 156.490 1.620 157.260 2.280 ;
        RECT 156.560 0.000 157.160 1.620 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 99.320 18.725 99.765 19.095 ;
        RECT 99.425 18.430 99.645 18.725 ;
        RECT 98.780 18.260 100.320 18.430 ;
      LAYER mcon ;
        RECT 99.435 18.805 99.630 19.030 ;
        RECT 98.860 18.260 100.240 18.430 ;
      LAYER met1 ;
        RECT 99.320 19.040 99.765 19.095 ;
        RECT 99.320 18.835 134.890 19.040 ;
        RECT 99.320 18.725 99.765 18.835 ;
        RECT 98.800 18.230 100.300 18.460 ;
        RECT 134.685 2.300 134.890 18.835 ;
        RECT 134.400 1.650 135.180 2.300 ;
      LAYER via ;
        RECT 134.600 1.800 135.010 2.190 ;
      LAYER met2 ;
        RECT 134.400 1.650 135.180 2.300 ;
      LAYER via2 ;
        RECT 134.600 1.800 135.010 2.190 ;
      LAYER met3 ;
        RECT 134.400 1.650 135.180 2.300 ;
      LAYER via3 ;
        RECT 134.600 1.800 135.010 2.190 ;
      LAYER met4 ;
        RECT 134.400 1.650 135.180 2.300 ;
        RECT 134.480 0.000 135.080 1.650 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.360000 ;
    PORT
      LAYER li1 ;
        RECT 85.080 22.180 85.735 22.575 ;
      LAYER mcon ;
        RECT 85.315 22.245 85.670 22.510 ;
      LAYER met1 ;
        RECT 85.080 22.180 85.735 22.575 ;
      LAYER via ;
        RECT 85.315 22.245 85.670 22.510 ;
      LAYER met2 ;
        RECT 85.080 22.180 85.735 22.575 ;
        RECT 85.210 14.970 85.450 22.180 ;
        RECT 85.210 14.730 112.920 14.970 ;
        RECT 112.680 3.300 112.920 14.730 ;
        RECT 112.400 2.720 113.000 3.300 ;
      LAYER via2 ;
        RECT 112.565 2.850 112.885 3.185 ;
      LAYER met3 ;
        RECT 112.400 2.720 113.000 3.300 ;
      LAYER via3 ;
        RECT 112.565 2.850 112.885 3.185 ;
      LAYER met4 ;
        RECT 112.400 0.000 113.000 3.300 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 85.960 22.055 88.000 22.225 ;
        RECT 85.980 21.320 87.980 22.055 ;
        RECT 90.110 21.680 91.650 21.850 ;
        RECT 85.990 15.710 87.980 21.320 ;
        RECT 90.125 20.720 91.630 21.680 ;
        RECT 98.775 21.670 99.615 21.840 ;
        RECT 101.225 21.730 102.765 21.900 ;
        RECT 99.110 21.015 99.280 21.670 ;
        RECT 90.180 15.710 91.540 20.720 ;
        RECT 99.040 20.665 99.385 21.015 ;
        RECT 101.245 20.900 102.745 21.730 ;
        RECT 95.000 17.775 96.540 17.945 ;
        RECT 95.020 16.950 96.520 17.775 ;
        RECT 95.030 15.710 96.515 16.950 ;
        RECT 101.250 15.710 102.740 20.900 ;
        RECT 85.190 12.955 86.980 14.105 ;
        RECT 85.395 11.670 86.810 12.955 ;
        RECT 85.395 10.255 103.735 11.670 ;
        RECT 102.320 9.495 103.735 10.255 ;
        RECT 101.815 8.085 103.975 9.495 ;
      LAYER mcon ;
        RECT 86.040 22.055 87.920 22.225 ;
        RECT 90.190 21.680 91.570 21.850 ;
        RECT 98.855 21.670 99.535 21.840 ;
        RECT 101.305 21.730 102.685 21.900 ;
        RECT 99.120 20.740 99.295 20.915 ;
        RECT 86.285 15.900 87.650 16.305 ;
        RECT 95.080 17.775 96.460 17.945 ;
        RECT 90.480 15.950 91.250 16.340 ;
        RECT 95.185 15.900 96.335 16.320 ;
        RECT 101.675 15.915 102.375 16.370 ;
        RECT 85.540 13.150 86.645 13.925 ;
        RECT 101.900 8.165 103.885 9.415 ;
      LAYER met1 ;
        RECT 85.980 22.025 87.980 22.255 ;
        RECT 90.130 21.650 91.630 21.880 ;
        RECT 98.795 21.640 99.595 21.870 ;
        RECT 101.245 21.700 102.745 21.930 ;
        RECT 99.040 20.665 99.385 21.015 ;
        RECT 99.095 20.480 99.335 20.665 ;
        RECT 97.830 20.240 99.335 20.480 ;
        RECT 95.020 17.745 96.520 17.975 ;
        RECT 51.640 16.490 52.685 16.715 ;
        RECT 97.830 16.490 98.070 20.240 ;
        RECT 51.640 15.710 102.750 16.490 ;
        RECT 51.640 15.475 52.685 15.710 ;
        RECT 85.190 12.955 86.980 15.710 ;
        RECT 101.840 8.135 103.945 9.445 ;
      LAYER via ;
        RECT 51.880 15.735 52.475 16.430 ;
        RECT 85.540 13.150 86.645 13.925 ;
      LAYER met2 ;
        RECT 51.640 15.475 52.685 16.715 ;
        RECT 85.190 12.955 86.980 14.105 ;
      LAYER via2 ;
        RECT 51.880 15.735 52.475 16.430 ;
        RECT 85.540 13.150 86.645 13.925 ;
      LAYER met3 ;
        RECT 51.640 15.475 52.685 16.715 ;
        RECT 57.210 13.665 84.070 31.440 ;
        RECT 85.280 13.665 86.980 14.105 ;
        RECT 57.210 13.250 86.980 13.665 ;
        RECT 57.210 11.040 84.070 13.250 ;
        RECT 85.280 12.955 86.980 13.250 ;
      LAYER via3 ;
        RECT 51.880 15.735 52.475 16.430 ;
        RECT 83.650 11.180 83.970 31.300 ;
      LAYER met4 ;
        RECT 49.000 16.490 50.500 220.760 ;
        RECT 51.640 16.490 52.685 16.715 ;
        RECT 49.000 15.705 52.685 16.490 ;
        RECT 49.000 5.000 50.500 15.705 ;
        RECT 51.640 15.475 52.685 15.705 ;
        RECT 83.570 11.100 84.050 31.380 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 100.185 24.375 100.515 24.440 ;
        RECT 100.810 24.375 101.020 24.380 ;
        RECT 100.185 24.205 101.020 24.375 ;
        RECT 85.330 23.940 88.610 24.110 ;
        RECT 100.185 24.100 100.515 24.205 ;
        RECT 86.045 23.345 87.925 23.940 ;
        RECT 88.890 23.530 89.225 23.805 ;
        RECT 88.950 23.345 89.165 23.530 ;
        RECT 86.045 23.160 89.165 23.345 ;
        RECT 86.045 22.695 87.925 23.160 ;
        RECT 100.810 22.810 101.020 24.205 ;
        RECT 85.960 22.525 88.000 22.695 ;
        RECT 100.140 22.640 101.020 22.810 ;
        RECT 98.285 21.820 98.600 22.155 ;
        RECT 94.100 21.450 97.380 21.620 ;
        RECT 95.000 21.170 96.380 21.450 ;
        RECT 95.000 20.995 97.205 21.170 ;
        RECT 95.000 20.730 96.380 20.995 ;
        RECT 94.950 20.560 96.490 20.730 ;
        RECT 97.035 20.630 97.205 20.995 ;
        RECT 97.035 20.440 97.210 20.630 ;
        RECT 94.950 20.090 96.490 20.260 ;
        RECT 94.970 19.285 96.470 20.090 ;
        RECT 97.040 20.070 97.210 20.440 ;
        RECT 98.355 20.070 98.535 21.820 ;
        RECT 100.140 20.070 100.370 22.640 ;
        RECT 100.810 22.270 101.020 22.640 ;
        RECT 100.670 21.870 101.040 22.270 ;
        RECT 97.040 19.900 100.370 20.070 ;
        RECT 95.115 18.985 96.330 19.285 ;
        RECT 95.115 18.975 97.735 18.985 ;
        RECT 95.115 18.805 97.740 18.975 ;
        RECT 95.115 18.415 96.330 18.805 ;
        RECT 95.000 18.245 96.540 18.415 ;
        RECT 97.535 17.320 97.740 18.805 ;
        RECT 98.355 18.305 98.545 19.900 ;
        RECT 98.755 19.895 100.175 19.900 ;
        RECT 98.325 17.925 98.600 18.305 ;
        RECT 98.780 17.790 100.320 17.960 ;
        RECT 98.795 17.320 100.305 17.790 ;
        RECT 97.535 17.135 100.305 17.320 ;
        RECT 98.795 16.950 100.305 17.135 ;
      LAYER mcon ;
        RECT 85.410 23.940 88.530 24.110 ;
        RECT 86.040 22.525 87.920 22.695 ;
        RECT 94.180 21.450 97.300 21.620 ;
        RECT 95.030 20.560 96.410 20.730 ;
        RECT 95.030 20.090 96.410 20.260 ;
        RECT 95.080 18.245 96.460 18.415 ;
        RECT 98.860 17.790 100.240 17.960 ;
      LAYER met1 ;
        RECT 85.350 23.910 88.590 24.140 ;
        RECT 85.980 22.495 87.980 22.725 ;
        RECT 94.120 21.420 97.360 21.650 ;
        RECT 94.970 20.530 96.470 20.760 ;
        RECT 94.970 20.060 96.470 20.290 ;
        RECT 95.020 18.215 96.520 18.445 ;
        RECT 98.800 17.760 100.300 17.990 ;
  END
END tt_um_lif
END LIBRARY

